library ieee;
use ieee.std_logic_1164.all;

package VGA_pkg is
   -- -------------------------------------------------------------------------
   -- Param�tres d'un �cran VGA de 640x480 � 60 Hz
   -- -------------------------------------------------------------------------
   
   -- La largeur de l'�cran, en pixels
   constant VGA_SCREEN_WIDTH : integer := 640;
   
   -- La hauteur de l'�cran, en pixels
   constant VGA_SCREEN_HEIGHT : integer := 480;
   
   -- Nombre de pixel sur l'�cran
   constant VGA_PIXEL_NUMBER : integer := VGA_SCREEN_WIDTH * VGA_SCREEN_HEIGHT;
   
   -- La valeur maximale de X, en pixels, rafra�chissement compris
   constant VGA_X_MAX : integer := 799;
   
   -- La valeur maximale de Y, en pixels, rafra�chissement compris
   constant VGA_Y_MAX : integer := 524;
   
   -- La coordonn�e X de d�but de l'impulsion de rafra�chissement horizontal
   constant VGA_HBL_START : integer := 659;
   
   -- La coordonn�e X de fin de l'impulsion de rafra�chissement horizontal
   constant VGA_HBL_END : integer := 755;

   -- La coordonn�e Y de d�but de l'impulsion de rafra�chissement vertical
   constant VGA_VBL_START : integer := 493;

   -- La coordonn�e Y de fin de l'impulsion de rafra�chissement vertical
   constant VGA_VBL_END : integer := 494;

   -- -------------------------------------------------------------------------
   -- D�finition des couleurs affichables
   -- -------------------------------------------------------------------------
   
   -- Type couleur
   --
   -- Cette structure fournit des champs pour les valeurs des composantes rouge, verte et bleue,
   -- et un champ indiquant si le pixel est opaque (visible) ou transparent (invisible).
   type VGAColor_t is record
      red : std_logic_vector(2 downto 0);
      green : std_logic_vector(2 downto 0);
      blue : std_logic_vector(1 downto 0);
      opaque : std_logic;
   end record VGAColor_t;

   -- D�finition de la couleur noire
   constant VGA_COLOR_BLACK : VGAColor_t := ("000", "000", "00", '1');

   -- D�finition de la couleur rouge
   constant VGA_COLOR_RED : VGAColor_t := ("111", "000", "00", '1');

   -- D�finition de la couleur verte
   constant VGA_COLOR_GREEN : VGAColor_t := ("000", "111", "00", '1');

   -- D�finition de la couleur bleue
   constant VGA_COLOR_BLUE : VGAColor_t := ("000", "000", "11", '1');

   -- D�finition de la couleur jaune
   constant VGA_COLOR_YELLOW : VGAColor_t := ("111", "111", "00", '1');

   -- D�finition de la couleur magenta
   constant VGA_COLOR_MAGENTA : VGAColor_t := ("111", "000", "11", '1');

   -- D�finition de la couleur cyan
   constant VGA_COLOR_CYAN : VGAColor_t := ("000", "111", "11", '1');

   -- D�finition de la couleur blanche
   constant VGA_COLOR_WHITE : VGAColor_t := ("111", "111", "11", '1');

   -- D�finition de la couleur "transparente"
   constant VGA_COLOR_TRANSPARENT : VGAColor_t := ("000", "000", "00", '0');
   
   -- -------------------------------------------------------------------------
   -- D�finition des caract�res affichables par VGATextPainter
   -- -------------------------------------------------------------------------
   
   -- Le nombre de caract�res diff�rents affichables
   constant VGA_CHARACTER_COUNT : integer := 128;
   
   -- La largeur d'un masque de caract�re, en points
   constant VGA_CHARACTER_WIDTH : integer := 5;
   
   -- La hauteur d'un masque de caract�re, en points
   constant VGA_CHARACTER_HEIGHT : integer := 7;

   -- La largeur d'affichage d'un caract�re � l'�cran, en points,
   -- pr�vue pour optimiser le taux d'occupation du FPGA.
   -- Cette largeur doit �tre une puissance de 2.
   constant VGA_CHARACTER_DISPLAY_WIDTH : integer := 8;

   -- La hauteur d'affichage d'un caract�re � l'�cran, en points,
   -- pr�vue pour optimiser le taux d'occupation du FPGA.
   -- Cette hauteur doit �tre une puissance de 2.
   constant VGA_CHARACTER_DISPLAY_HEIGHT : integer := 8;
	
	
	-- d�claration type : tableau d'entier et de couleur ( 16 indice ) 
	type int_array is array(0 to 15) of integer;
	
	type color_array is array (0 to 15) of VGAColor_t;	
	
	type full_screen_array_t is array (0 to VGA_PIXEL_NUMBER-1) of VGAColor_t;	

   type VGAString_t is array (integer range <>) of integer range 0 to VGA_CHARACTER_HEIGHT * VGA_CHARACTER_COUNT - 1;
  
   type VGACharacterBitmap_t is array(0 to VGA_CHARACTER_HEIGHT * VGA_CHARACTER_COUNT - 1)
      of std_logic_vector(0 to VGA_CHARACTER_WIDTH - 1);
   
   constant VGA_CHARACTER_BITMAP : VGACharacterBitmap_t := (
      -- Caract�re 0 : ' '
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 1 (129) : '�'
      "10001", -- *   *
      "00000", -- 
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10011", -- *  **
      "01101", --  ** *

      -- Caract�re 2 (130) : '�'
      "00010", --    *
      "00100", --   *
      "01110", --  ***
      "10001", -- *   *
      "11111", -- *****
      "10000", -- *   
      "01110", --  ***
      
      -- Caract�re 3 (131): '�'
      "01110", --  ***
      "00000", -- 
      "01110", --  ***
      "00001", --     *
      "01111", --  ****
      "10001", -- *   *
      "01111", --  ****

      -- Caract�re 4 (132): '�'
      "01010", --  * *
      "00000", -- 
      "01110", --  ***
      "00001", --     *
      "01111", --  ****
      "10001", -- *   *
      "01111", --  ****

      -- Caract�re 5 (133): '�'
      "01000", --  *
      "00100", --   *
      "01110", --  ***
      "00001", --     *
      "01111", --  ****
      "10001", -- *   *
      "01111", --  ****

      -- Caract�re 6 (134): ''
      "00100", --   *
      "00000", -- 
      "01110", --  ***
      "00001", --     *
      "01111", --  ****
      "10001", -- *   *
      "01111", --  ****

      -- Caract�re 7 (135) : '�'
      "00000", -- 
      "00000", -- 
      "01110", --  ***
      "10000", -- *   
      "10001", -- *   *
      "01110", --  ***
      "11000", -- ** 

      -- Caract�re 8 (136) : '�'
      "01110", --  ***
      "00000", -- 
      "01110", --  ***
      "10001", -- *   *
      "11111", -- *****
      "10000", -- *   
      "01110", --  ***

      -- Caract�re 9 (137) : '�'
      "01010", --  * *
      "00000", -- 
      "01110", --  ***
      "10001", -- *   *
      "11111", -- *****
      "10000", -- *   
      "01110", --  ***

      -- Caract�re 10 (138) : '�'
      "01000", --  *
      "00100", --   *
      "01110", --  ***
      "10001", -- *   *
      "11111", -- *****
      "10000", -- *   
      "01110", --  ***

      -- Caract�re 11 (139): '�'
      "01010", --  * *
      "00000", -- 
      "01100", --  **
      "00100", --   * 
      "00100", --   *
      "00100", --   *
      "01110", --  ***

      -- Caract�re 12 (140) : '�'
      "01110", --  ***
      "00000", -- 
      "01100", --  **
      "00100", --   * 
      "00100", --   *
      "00100", --   *
      "01110", --  ***

      -- Caract�re 13 : Fl�che haut
      "00100", --   *
      "01110", --  ***
      "10101", -- * * *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      
      -- Caract�re 14 : Fl�che bas
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "10101", -- * * *
      "01110", --  ***
      "00100", --   *
            
      -- Caract�re 15 : Fl�che droite
      "00000", -- 
      "00100", --   *
      "00010", --    *
      "11111", -- *****
      "00010", --    *
      "00100", --   *
      "00000", -- 
      
      -- Caract�re 16 : Fl�che gauche
      "00000", -- 
      "00100", --   *
      "01000", --  *
      "11111", -- *****
      "01000", --  *
      "00100", --   *
      "00000", -- 

      -- Caract�re 17 : Croix de multiplication
      "00000", -- 
      "10001", -- *   *
      "01010", --  * *
      "00100", --   *
      "01010", --  * *
      "10001", -- *   *
      "00000", -- 
      
      -- Caract�re 18 : Division
      "00000", -- 
      "00100", --   * 
      "00000", -- 
      "11111", -- *****
      "00000", -- 
      "00100", --   *
      "00000", -- 

      -- Caract�re 19 (147) : '�'
      "01110", --  ***
      "00000", -- 
      "01110", --  ***
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***

      -- Caract�re 20 (148) : '�'
      "01010", --  * *
      "00000", -- 
      "01110", --  ***
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***
      
      -- Caract�re 21 : Diamant
      "00000", -- 
      "00100", --   *
      "01010", --  * *
      "10001", -- *   *
      "01010", --  * *
      "00100", --   *
      "00000", -- 

      -- Caract�re 22 (150) : '�'
      "01110", --  ***
      "00000", -- 
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10011", -- *  **
      "01101", --  ** *

      -- Caract�re 23 (151) : '�'
      "01000", --  *
      "00100", --   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10011", -- *  **
      "01101", --  ** *
           
      -- Caract�re 24 : Grand rectangle
      "11111", -- *****
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "11111", -- *****
      
      -- Caract�re 25 : Petit rectangle
      "00000", -- 
      "01110", --  ***
      "01010", --  * *
      "01010", --  * *
      "01010", --  * *
      "01110", --  ***
      "00000", -- 
      
      -- Caract�re 26 : Grand carr�
      "00000", -- 
      "11111", -- *****
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "11111", -- *****
      "00000", -- 
      
      -- Caract�re 27 : Petit carr�
      "00000", -- 
      "00000", -- 
      "01110", --  ***
      "01010", --  * *
      "01110", --  ***
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 28 : Point central
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00100", --   * 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 29 : Sup�rieur ou �gal (non ASCII)
      "10000", -- *
      "01000", --  *
      "00100", --   *
      "00010", --    *
      "11111", -- *****
      "00000", -- 
      "11111", -- *****
      
      -- Caract�re 30 : Inf�rieur ou �gal (non ASCII)
      "00001", --     *
      "00010", --    *
      "00100", --   *
      "01000", --  *
      "11111", -- *****
      "00000", -- 
      "11111", -- *****
      
      -- Caract�re 31 : Diff�rent
      "00000", -- 
      "00000", -- 
      "00010", --    *
      "11111", -- *****
      "00100", --   *
      "11111", -- *****
      "01000", --  *
      
      -- Caract�re 32 : ' '
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 

      -- Caract�re 33 : '!'
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00000", -- 
      "00100", --   *
      
      -- Caract�re 34 : '"'
      "01010", --  * *
      "01010", --  * *
      "01010", --  * *
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 35 : '#'
      "01010", --  * *
      "01010", --  * *
      "11111", -- *****
      "01010", --  * *
      "11111", -- *****
      "01010", --  * *
      "01010", --  * *
      
      -- Caract�re 36 : '$'
      "00100", --   *
      "01110", --  ****
      "10100", -- * * 
      "01110", --  ***
      "00101", --   * *
      "11110", -- ****
      "00100", --   *
      
      -- Caract�re 37 : '%'
      "11000", -- **
      "11001", -- **  *
      "00010", --    *
      "00100", --   *
      "01000", --  *
      "10011", -- *  **
      "00011", --    **
      
      -- Caract�re 38 : '&'
      "01100", --  **
      "10010", -- *  *
      "10100", -- * *
      "01000", --  *
      "10101", -- * * *
      "10010", -- *  *
      "01101", --  ** *
      
      -- Caract�re 39 : '''
      "01100", -- **
      "00100", --  *
      "01000", -- *
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 40 : '('
      "00010", --    *
      "00100", --   *
      "01000", --  *
      "01000", --  *
      "01000", --  *
      "00100", --   *
      "00010", --    *
      
      -- Caract�re 41 : ')'
      "01000", --  *
      "00100", --   *
      "00010", --    *
      "00010", --    *
      "00010", --    *
      "00100", --   *
      "01000", --  *
      
      -- Caract�re 42 : '*'
      "00000", -- 
      "00100", --   *
      "10101", -- * * *
      "01110", --  *** 
      "10101", -- * * *
      "00100", --   *
      "00000", -- 
      
      -- Caract�re 43 : '+'
      "00000", -- 
      "00100", --   *
      "00100", --   * 
      "11111", -- *****
      "00100", --   * 
      "00100", --   *
      "00000", -- 
      
      -- Caract�re 44 : ','
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "01100", -- **
      "00100", --  *
      "01000", -- *
      
      -- Caract�re 45 : '-'
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "11111", -- *****
      "00000", -- 
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 46 : '.'
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", --
      "01100", --  **
      "01100", --  **
      "00000", --
      
      -- Caract�re 47 : '/'
      "00000", -- 
      "00001", --     *
      "00010", --    *
      "00100", --   *
      "01000", --  *
      "10000", -- *
      "00000", -- 

      -- Caract�re 48 : '0'
      "01110", --  ***
      "10001", -- *   *
      "10011", -- *  **
      "10101", -- * * *
      "11001", -- **  *
      "10001", -- *   *
      "01110", --  ***
      
      -- Caract�re 49 : '1'
      "00100", --   * 
      "01100", --  **
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "01110", --  ***
      
      -- Caract�re 50 : '2'
      "01110", --  ***
      "10001", -- *   *
      "00001", --     *
      "00010", --   *
      "00100", --  *
      "01000", -- *
      "11111", -- *****
      
      -- Caract�re 51 : '3'
      "11111", -- *****
      "00010", --    *
      "00100", --   *
      "00010", --    *
      "00001", --     *
      "10001", -- *   *
      "01110", --  ***
      
      -- Caract�re 52 : '4'
      "00010", --    * 
      "00110", --   **
      "01010", --  * *
      "10010", -- *  *
      "11111", -- *****
      "00010", --    *
      "00010", --    *
      
      -- Caract�re 53 : '5'
      "11111", -- *****
      "10000", -- *
      "11110", -- ****
      "00001", --     *
      "00001", --     *
      "10001", -- *   *
      "01110", --  ***
      
      -- Caract�re 54 : '6'
      "00110", --   **
      "01000", --  *
      "10000", -- *
      "11110", -- ****
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***
      
      -- Caract�re 55 : '7'
      "00110", -- *****
      "01000", --     *
      "10000", --    *
      "11110", --   *
      "10001", --  *
      "10001", -- *
      "01110", -- *
      
      -- Caract�re 56 : '8'
      "01110", --  *** 
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***
      
      -- Caract�re 57 : '9'
      "01110", --  *** 
      "10001", -- *   *
      "10001", -- *   *
      "01111", --  ****
      "00001", --     *
      "00010", --    *
      "01100", --  **
      
      -- Caract�re 58 : ':'
      "00000", -- 
      "01100", --  **
      "01100", --  **
      "00000", --
      "01100", --  **
      "01100", --  **
      "00000", --
      
      -- Caract�re 59 : ';'
      "00000", -- 
      "01100", --  **
      "01100", --  **
      "00000", --
      "01100", --  **
      "00100", --   *
      "01000", --  *

      -- Caract�re 60 : '<'
      "00010", --    *
      "00100", --   *
      "01000", --  *
      "10000", -- *
      "01000", --  *
      "00100", --   *
      "00010", --    *

      -- Caract�re 61 : '='
      "00000", -- 
      "00000", -- 
      "11111", -- *****
      "00000", -- 
      "11111", -- *****
      "00000", -- 
      "00000", -- 

      -- Caract�re 62 : '>'
      "01000", --  *
      "00100", --   *
      "00010", --    *
      "00001", --     *
      "00010", --    *
      "00100", --  *
      "01000", -- *

      -- Caract�re 63 : '?'
      "01110", --  ***
      "10001", -- *   *
      "00001", --     *
      "00010", --    *
      "00100", --   *
      "00000", -- 
      "00100", --   *

      -- Caract�re 64 : '@'
      "01110", --  ***
      "10001", -- *   *
      "00001", --     *
      "01101", --  ** *
      "10101", -- * * *
      "10101", -- * * *
      "01110", --  ***

      -- Caract�re 65 : 'A'
      "01110", --  ***
      "10001", -- *   *
      "10001", -- *   *
      "11111", -- *****
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *

      -- Caract�re 66 : 'B'
      "11110", -- ****
      "10001", -- *   *
      "10001", -- *   *
      "11110", -- ****
      "10001", -- *   *
      "10001", -- *   *
      "11110", -- ****

      -- Caract�re 67 : 'C'
      "01110", --  ***
      "10001", -- *   *
      "10000", -- *
      "10000", -- *
      "10000", -- *
      "10001", -- *   *
      "01110", --  ***

      -- Caract�re 68 : 'D'
      "11110", -- ****
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "11110", -- ****

      -- Caract�re 69 : 'E'
      "11111", -- *****
      "10000", -- *
      "10000", -- *
      "11110", -- ****
      "10000", -- *
      "10000", -- *
      "11111", -- *****

      -- Caract�re 70 : 'F'
      "11111", -- *****
      "10000", -- *
      "10000", -- *
      "11110", -- ****
      "10000", -- *
      "10000", -- *
      "10000", -- *

      -- Caract�re 71 : 'G'
      "01110", --  ***
      "10001", -- *   *
      "10000", -- *
      "10111", -- * ***
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***

      -- Caract�re 72 : 'H'
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "11111", -- *****
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *

      -- Caract�re 73 : 'I'
      "01110", --  *** 
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "01110", --  ***

      -- Caract�re 74 : 'J'
      "00111", --   ***
      "00010", --    *
      "00010", --    *
      "00010", --    *
      "00010", --    *
      "10010", -- *  *
      "01100", --  ** 

      -- Caract�re 75 : 'K'
      "10001", -- *   *
      "10010", -- *  *
      "10100", -- * *
      "11000", -- **
      "10100", -- * *
      "10010", -- *  *
      "10001", -- *   *

      -- Caract�re 76 : 'L'
      "10000", -- *
      "10000", -- *
      "10000", -- *
      "10000", -- *
      "10000", -- *
      "10000", -- *
      "11111", -- *****

      -- Caract�re 77 : 'M'
      "10001", -- *   *
      "11011", -- ** **
      "10101", -- * * *
      "10101", -- * * *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *

      -- Caract�re 78 : 'N'
      "10001", -- *   *
      "10001", -- *   *
      "11001", -- **  *
      "10101", -- * * *
      "10011", -- *  **
      "10001", -- *   *
      "10001", -- *   *

      -- Caract�re 79 : 'O'
      "01110", --  ***
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***

      -- Caract�re 80 : 'P'
      "11110", -- ****
      "10001", -- *   *
      "10001", -- *   *
      "11110", -- ****
      "10000", -- *
      "10000", -- *
      "10000", -- *

      -- Caract�re 81 : 'Q'
      "01110", --  ***
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10101", -- * * *
      "10010", -- *  * 
      "01101", --  ** *

      -- Caract�re 82 : 'R'
      "11110", -- ****
      "10001", -- *   *
      "10001", -- *   *
      "11110", -- ****
      "10100", -- * *
      "10010", -- *  *
      "10001", -- *   *

      -- Caract�re 83 : 'S'
      "01110", --  ***
      "10001", -- *   *
      "10000", -- *
      "01110", --  *** 
      "00001", --     *
      "10001", -- *   *
      "01110", --  ***

      -- Caract�re 84 : 'T'
      "11111", -- *****
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *

      -- Caract�re 85 : 'U'
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***

      -- Caract�re 86 : 'V'
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "01010", --  * * 
      "00100", --   *

      -- Caract�re 87 : 'W'
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10101", -- * * *
      "10101", -- * * *
      "11011", -- ** **
      "10001", -- *   *

      -- Caract�re 88 : 'X'
      "10001", -- *   *
      "10001", -- *   *
      "01010", --  * *
      "00100", --   *
      "01010", --  * *
      "10001", -- *   *
      "10001", -- *   *

      -- Caract�re 89 : 'Y'
      "10001", -- *   *
      "10001", -- *   *
      "01010", --  * *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *

      -- Caract�re 90 : 'Z'
      "11111", -- *****
      "00001", --     *
      "00010", --    *
      "00100", --   *
      "01000", --  *
      "10000", -- *
      "11111", -- *****

      -- Caract�re 91 : '['
      "01110", --  ***
      "01000", --  *
      "01000", --  *
      "01000", --  *
      "01000", --  *
      "01000", --  *
      "01110", --  ***

      -- Caract�re 92 : '\'
      "00000", -- 
      "10000", -- *
      "01000", --  *
      "00100", --   *
      "00010", --    *
      "00001", --     *
      "00000", -- 

      -- Caract�re 93 : ']'
      "01110", --  ***
      "00010", --    *
      "00010", --    *
      "00010", --    *
      "00010", --    *
      "00010", --    *
      "01110", --  ***

      -- Caract�re 94 : '^'
      "00100", --   *
      "01010", --  * *
      "10001", -- *   *
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 95 : '_'
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "11111", -- *****
      
      -- Caract�re 96 : '`'
      "00110", --  **
      "00100", --  *
      "00010", --   *
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "00000", -- 
      
      -- Caract�re 97 : 'a'
      "00000", -- 
      "00000", -- 
      "01110", --  ***
      "00001", --     *
      "01111", --  ****
      "10001", -- *   *
      "01111", --  ****

      -- Caract�re 98 : 'b'
      "10000", -- *
      "10000", -- *
      "10110", -- * **
      "11001", -- **  *
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  *** 

      -- Caract�re 99 : 'c'
      "00000", -- 
      "00000", -- 
      "01110", --  ***
      "10000", -- *   
      "10000", -- *
      "10001", -- *   *
      "01110", --  *** 

      -- Caract�re 100 : 'd'
      "00001", --     *
      "00001", --     *
      "01101", --  ** *
      "10011", -- *  **
      "10001", -- *   *
      "10001", -- *   *
      "01111", --  **** 
      
      -- Caract�re 101 : 'e'
      "00000", -- 
      "00000", -- 
      "01110", --  ***
      "10001", -- *   *
      "11111", -- *****
      "10000", -- *   
      "01110", --  ***

      -- Caract�re 102 : 'f'
      "00010", --    *
      "00101", --   * *
      "00100", --   *
      "01110", --  ***
      "00100", --   *
      "00100", --   *
      "00100", --   *
      
      -- Caract�re 103 : 'g'
      "00000", -- 
      "00000", -- 
      "01111", --  ****
      "10001", -- *   *
      "01111", --  ****
      "00001", --     *
      "01110", --  ***

      -- Caract�re 104 : 'h'
      "10000", -- *
      "10000", -- *
      "10110", -- * **
      "11001", -- **  *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *

      -- Caract�re 105 : 'i'
      "00100", --   *
      "00000", -- 
      "01100", --  **
      "00100", --   * 
      "00100", --   *
      "00100", --   *
      "01110", --  ***
      
      -- Caract�re 106 : 'j'
      "00010", --    * 
      "00000", -- 
      "00010", --    * 
      "00010", --    *
      "00010", --    *
      "10010", -- *  *
      "01100", --  **

      -- Caract�re 107 : 'k'
      "10000", -- *
      "10000", -- *
      "10010", -- *  *
      "10100", -- * *
      "11000", -- **
      "10100", -- * *
      "10010", -- *  *

      -- Caract�re 108 : 'l'
      "01100", --  **
      "00100", --   *
      "00100", --   *
      "00100", --   * 
      "00100", --   *
      "00100", --   *
      "01110", --  ***

      -- Caract�re 109 : 'm'
      "00000", -- 
      "00000", -- 
      "11010", -- ** *
      "10101", -- * * *
      "10101", -- * * *
      "10101", -- * * *
      "10101", -- * * *

      -- Caract�re 110 : 'n'
      "00000", -- 
      "00000", -- 
      "10110", -- * **
      "11001", -- **  *
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *

      -- Caract�re 111 : 'o'
      "00000", -- 
      "00000", -- 
      "01110", --  ***
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "01110", --  ***

      -- Caract�re 112 : 'p'
      "00000", -- 
      "00000", -- 
      "11110", -- ****
      "10001", -- *   *
      "11110", -- ****
      "10000", -- *   
      "10000", -- *

      -- Caract�re 113 : 'q'
      "00000", -- 
      "00000", -- 
      "01111", --  ****
      "10001", -- *   *
      "01111", --  ****
      "00001", --     *   
      "00001", --     *

      -- Caract�re 114 : 'r'
      "00000", -- 
      "00000", -- 
      "01011", --  * **
      "01100", --  **
      "01000", --  *
      "01000", --  *
      "01000", --  *
      
      -- Caract�re 115 : 's'
      "00000", -- 
      "00000", -- 
      "01111", --  ****
      "10000", -- *
      "01110", --  ***
      "00001", --     *
      "11110", -- ****

      -- Caract�re 116 : 't'
      "00000", -- 
      "00100", --   *
      "01110", --  ***
      "00100", --   * 
      "00100", --   *
      "00101", --   * *
      "00010", --    *

      -- Caract�re 117 : 'u'
      "00000", -- 
      "00000", -- 
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "10011", -- *  **
      "01101", --  ** *

      -- Caract�re 118 : 'v'
      "00000", -- 
      "00000", -- 
      "10001", -- *   *
      "10001", -- *   *
      "10001", -- *   *
      "01010", --  * *
      "00100", --   *

      -- Caract�re 119 : 'w'
      "00000", -- 
      "00000", -- 
      "10001", -- *   *
      "10001", -- *   *
      "10101", -- * * *
      "10101", -- * * *
      "01010", --  * *

      -- Caract�re 120 : 'x'
      "00000", -- 
      "00000", -- 
      "11001", -- **  *
      "00110", --   ** 
      "00100", --   *
      "01100", --  **
      "10011", -- *  **

      -- Caract�re 121 : 'y'
      "00000", -- 
      "00000", -- 
      "10001", -- *   *
      "01001", --  *  *
      "00110", --   **
      "00100", --   *
      "11000", -- **

      -- Caract�re 122 : 'z'
      "00000", -- 
      "00000", -- 
      "11111", -- *****
      "00010", --    * 
      "00100", --   *
      "01000", --  * 
      "11111", -- *****

      -- Caract�re 123 : '{'
      "00011", --    **
      "00100", --   *
      "00100", --   *
      "11000", -- **
      "00100", --   *
      "00100", --   *
      "00011", --    **

      -- Caract�re 124 : '|'
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *
      "00100", --   *

      -- Caract�re 125 : '}'
      "11000", -- **
      "00100", --   *
      "00100", --   *
      "00011", --    **
      "00100", --   *
      "00100", --   *
      "11000", -- **

      -- Caract�re 126 : '~'
      "00000", -- 
      "00000", -- 
      "00000", -- 
      "01010", --  * * 
      "10100", -- * *
      "00000", --
      "00000", --

      -- Caract�re 127 : DEL
      "11111", -- ***** 
      "11111", -- ***** 
      "11111", -- ***** 
      "11111", -- ***** 
      "11111", -- ***** 
      "11111", -- ***** 
      "11111"  -- ***** 
   );
end VGA_pkg;

